

module Plain_Text(


    );
endmodule